module vna

fn unit<T>() {}
