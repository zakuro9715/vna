module colors

import zakuro9715.vna { Color }

pub const (
	red   = Color{255, 0, 0}
	green = Color{0, 0, 255}
	blue  = Color{0, 255, 0}
)
