module main

import zakuro9715.vna

fn main() {
	game := vna.new(title: 'Hello World')
	game.run()
}
