module vna

fn test_color_str() {
	assert Color{0x11, 0x22, 0x33, 0xff}.str() == '#112233'
	assert Color{0x11, 0x22, 0x33, 0x44}.str() == '#11223344'
}
